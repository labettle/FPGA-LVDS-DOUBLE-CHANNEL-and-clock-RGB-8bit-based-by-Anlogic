module idelay_ctrl (
    input wire    I_clk,
    input wire    I_rst,

    input wire    I_dpa_start,
    input wire    I_lane_match,
    output reg    O_lane_dpa_done,
    
    output wire[7:0]	O_idelay_num,
    output wire	[7:0]	O_eye_taps
);
	
    
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Anlogic"
`pragma protect encrypt_agent_info = "Anlogic Encryption Tool anlogic_2019"
`pragma protect key_keyowner = "Anlogic", key_keyname = "anlogic-rsa-001"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`pragma protect key_block
LmbsqOWpj/6BLMfk860QqCFL+t4wq87o+nLgXnzADKMSNReTfysyXTofH5eKUFTs
1r6elHg+4BFFbdXGxASwgJ77mKLU1cks0oSrq/YnHvXrc24wxXM2Or1HGBieo8Oy
gWojI/xJXiKDl+caloCIQAUH8dsU98CjEDFUryYnJog=
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "CDS_RSA_KEY_VER_1"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 256)
`pragma protect key_block
nhEWjk88fw9wj+NkOZbtfm6B5js+mmgpljANmMSmX0aALxQzsWUHUkwjWAN1q3bG
SxPxz5eDC2CDd0M/Uz351jZh1WbLkMp+LUE7GKGHSoEtn3MMwcrHMmPt070DI6Me
qib5ZJ/8Pv3/Hi0+G1tgNE+TssZvgYl4naXXOfe0Ue6iqzjioIHCMneXJNda2uPg
LaG1RB+mm7bwev+xVl3Ptos8ymeNkL6XddeCPfJyeBUoJ+ByBejjmoSu6ohyJyBj
ZKDgze5PRvGmRlHwMF+j26pSFoEWS3JB/x3OYihcceCT7SzJ9rhd34FxFYWtyfwY
HoHf0dadQQNgHTJfoDzKiQ==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`pragma protect key_block
KzWPiDNobtRxHUv3G4ZvNrzjGW6ePyrfoEl3EqkdEL2EfHJ7unAozUHfMkrpCTgA
2N5uW7w/BWuMJhFCVQoDShTnlBuwYIP6NZicZag6m+Zo5IsAGGJivLaPg85yHI8c
JjJJXrtfpVnWlw0F9ITX2dKF3qkPkB4ZlflKNINFo+M=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 256)
`pragma protect key_block
AgdWUXdNPHaS96mKIkvOUVIfCqKjXYKesux5R6oJXT5gAqWvp3ABQlwwxbg3Rodx
WLlch8+ZMAqMGrNBu7RJwje9PQWQoJEcR2JftqOwUx8D8jZZpQXM5gE5amoOA18n
QwLluBEP+UmRsx+z6S8UBssTcrbbk0B0Spk0aSCQ/q7ZtCbPBWGs/+7BAOfqfRME
IXr4RyJO7qREVoyRhEEzcgnN5cHs72dFPgrp5VCPCygut65EMogx+2jbOfb3UFQT
le3xLgSzCK9EHL4UJGL5iLxPe33cuT9GUKi6XT/FMjY93WLYVkqvdt0pRtRDpxdG
vdKZBqrN23sZspddZ5vdEA==
`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`pragma protect key_block
qgsRFlmd/on2iTEzprt3f+oOVGAkwUX3qCjqoJVykI5/3vH8oVWXnQTsnbUo5KMW
RyGgY3g9c01qd17CoLqcZtXmUQXqmTq4nEaQqzG+ZmjuF3OaS4bAiVoiWpcst/5D
fmNL3viinrYgOAJ+//49OTFhlncpIpM9x2DJ1542ZNU=
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 9840)
`pragma protect data_block
FWhvO1XClkmQKqufO9Yb45+kUlAenBlkwjncJQqyX7kaWiart0vGlvZGu1dHAWNC
zzbSFzoQ3uS4H8FfxcdzDW2Q62nbD9aiRCD+eWw70w9v7FVHLGw9nOWQ2Kg/4SWr
6YjMaFJdyo7JcvFdkRjPepMP6D9XlkTmQyTXpU/r7yLqTTmkQqdO2HEO3DGOAQtf
Eg7qUNcFFJhlRfJ2tfNuU/nwzU4ouxTjCdN2TJSiiUmo/HDs6gBTApUPPcbWatDX
LMFaCz2134Knul3rIU253KRAM0czwXa+uypM1L98FwgNe4WrA8C0W4lamPTYQ1Nn
8sHl3NebFlMDTXnVq4ETArkhJs2G3/OD51oqLdH6CiH/tSM2pXHTBZ2hSVsUaOJq
R9Lf+/Xi4R8tEsg6xerG3mkjzPWBT0RextbdbqYkzDhz4dp845YJ1IMPLukQXxPs
op+HZOapEGVL/OLLwpfeesOMd3iypxVVmk4R43ZHojfvD98KNd1auT/xG/u+ZK5D
F1WXWERl0PbWTao7y+S/dJzeafeuRNfokv+8Y2Q4Le8DkEZr6wBzKmtEwEYVX+3j
5oBDu4s0vE+a7ISXNTJdJT4O10mW6XSiizQRJt+i8xcetd9lh96+W+CDYVJueMui
LqtyqArQDuZ/eJ2H+pR4+h1DzN1UpPwjkF/ClINoA+g3jh3yBDr4MuYzW7EslXdj
yym/7iGTMdH+RZUwkmEPF7Q8AgYF+HQcHJCtLU9s02ghgKBBkPnynMKWWeO44BCy
4wgQE2A1fPz73XnG+BPKlcj9fzE9C7K2urRh5UMYNiTaqrmqJOYnTz8ZGpl29Kzb
o7iE1aNHrxcUiqKxr8o0pkVfEHdSSFD0Ljg99eWVOMmTUcRp4LkFajaU8yanDk6D
76OsLK+8HATL1IrK0A5UZEpVshLhEJqSatEMA0WxWB2oAHBESnA0d9o9uActxwfQ
QSKiJrhAk8A3SCDy9EqXK3GSk3u11OHshVbOJwl2Qg4f5o/rYwR+KK7XG5maovjJ
2oTAoBOHAmqIO5ezxb5STnQ794CtmtqjtKG3gPkbukwJ9Kad1mi02p9U7R7MBX9u
l9oZUZAt3teKQDAJoC5ECOA6laejru1HGiyrH4IQ1jYrOmaEd8yOfsKhrsVrgHoR
T9yVDRPqhbEkZtE6Pbqdr6+vcS1iUxD8JD6sKaJKFiT4M51AT1GWbXnoPEFXfFIa
ggU4JE4DNA5cWX5v6+omdRWl9F0mTisu4xMZdKx+wmjoA6/9lNyHtugGH/NiIGcN
77Gk2bjzlP3ZqwvPIWLmc8syVWoTKBqb7VkoEZ4OVlZUzIY0cN7UJlX6BdVDrSKR
Ihbxu63oL3BJBVaffPMLtk7n+2ehdaP/Jw8xWCWVFqyTaX/5aZ1AGEhPYYU8awBv
k68IyYcU0Ae+B0WJcNfjlvmiDlSLIpHYHHjx1J7CAlU66wgc+7sv952JzsZ9/kx0
F/OqJ6IBiNB5Dm5XXIg6lui64ofOS+IViBNij21H9M3IZzVzL0PzmRfILdHWs/Ey
FV9j9g63VkIYWlGrXNQa9E+3H8boxIa4if6/LLuXNiP3X+Bur74fdweCcVKOZCVj
JqBJZ5hpAGK9KPJLz7xkzl7Q/hRpHOUvFR5X84OeM3ChT9ExiBj6wBjL5OxZqAze
B+kzjO/vBCPJ0XhoDRnvJFBRcBnj7VH2x1stqehQVMzernTt8Ekz56oLp75bbDk0
E2Qx6h+qRIjWnSPsuDzl2v4eXt9438yUiV4VKN5kqCmyJfvAfxYUFfKPOcapda7g
QywISsG9Yz2oDLGZGvrKVMx2RSpS9FcE7xJhdcA2HzPn+hs3W+rZ2bAKpww91IUD
2ObuBoPCDCb7HlG6Lux01WBxpoRIgS0VEjgt9PEJHn5pXjLxlEW8U5BeUnkTMR4g
V400yFF6gJvW3Bcj1nvzB+A21uluoQWj7K2uXrVQscPyZqR4twyycECAPBjMcdNM
ZFbr6LPgs9MjRn1XMn+RnhEm2ekA8qmrhIplP/nKfCTO2xP6aZomXlRXrQOfsGLY
BR1OkXv1RLzVwMfLzRjY6+95JydqcC3ocERJxXOU5x5VIMbCyZUWCs69GrnwAmVn
L+8NxTiY4sJsYFX5m6mlxILGruvc71yUo5VLCze/7BPmAnqV/06p6tpX7+qgM2yS
NzlQVB5C7Lku94/SwAAozdPJLG5x6QeKJ0YCDS1MO5S2g9nxTXz1lp7YIIFt4PGH
CDC0cpCfmZo4IrBnq7feBHng5HgAJj5PBSY5W75PpNWYV3v9LhBOjQWHqlp9F/el
6NAm7EE0pIZh4jTDGCJ2mc+lFQCbqryQMhNa+2ACmtZnpTLIEDMO56aBhrNPVGsm
QYs6rMYXcSzoGrpABjtJJcygH4e/ordITUiIb67ROHzzpnxKlugYL79dyy/+oEDR
uR5pz6kksm8rGg+VIu8zeZ//PYOFESImidn4LCHtZs8Egl5Ss/Z9xmfNjF2hHnyO
4oYJ/fBVzjkLzujrOULHDi0Ku1Epk/WdHH3RkbXU/CprBwHrg7Si6cX2Frb4KrFb
CByn7ZcvtZAyPirPYCk/S0+3N9Zw5CWAUYqRoFsrZZprzvrkFx+eydKmUG+XvFR6
YwD2Ngw2cTApTEhbfBw+xffV3yC8QsfIOXFfPNGIETLs8SvxFbVt6JqVq+x+yNZ6
wQcPF67ulcU1j1h7dlAkjRdDe1Y1w7OH99CFLEP+gRK0NjtKy5YROccPN32NmwVo
Ezg0upnK3VK/WjK0r6ixooDNlm/3jXaUTQi3T9xg9aiqMZEsVs3LfiDhNciyLHkG
HccOP3tF7TStb/JGWDtYgZs/0dAkjPWyewCx6OIvD7GykQvVDF6005RpbwchlU8W
zHKxFxYbhjIf/uw8Tfr8ADe6Sh0jBIIfOa7Q/Cm2I10uiZ2DIdIEHV/Frgcm4PVi
PqdSBfOTScG4+6NPIhRWy7PiMnHCXRm6vJ3tD4ivULQlNox/nS70WvguyAm0Sb9D
Jj/dwzV/vDsiU6kK2YHj8IPGoax2Bftpj1RbwSesLiP4vefCXeshWatc/l0FOS7B
4pDANfpvFb0uBmp/+qc2eorJOi2UcsvyVkz2i/+S/50HlWcr5GJl5hsf5yAdamKm
FLx5Eh81D6w81BzxPYVKaDM8A56EIynHsSIwA50t5Ft3TWIf/lOWMA+BMPHccLwT
Myx3Oqn7Atcm01KvqkMIDEPckjWY9rpC3peB4f/hiXZAIhq8iQHseufEi5dR/YrW
1haqNcUPIGjXX3/jfDjy1SmpiGdUAesvsLcpj9/0d21oAFZIIx4KrOQ/diiE7vDd
S5nIkytghGAVqnA26Jw+Bzb6fT/G9OnbBTa3vv5A7Pzv/b74TUlHdIKi9tPyWm7n
/YT/vC6mbaBhEkPTQlZa4NmqkN1f2nk2WU9BaJv230SF/Wxl49Oy2KfSid8pod+P
Thdx5+IKpRcxbgoLLvilnnSup1/ixmePT5uOseLmzhJyv3jHLQjgHlufF7LcAObG
40bwq1q0G8VgvmCTt9TYD6HeFZrEuNSGsLbQmu7tpOpMZsS7+UCoc+VhFU3qU9Mk
/sqhvABPMh32q/hEOfTFz+C9rC0YkAdB/GpAd3Hkz3cTXnSZ1ZiQ0OK7ESQX9f2d
jH+2CW5p3E86AFXNKHnnTuUvDu5eAceWfNY/9KoG91zZI8jmSmajdAlX5WjPgS+1
oPzsJq3DIlRmLC5BAzLFVhD9g6KwRux5VuFNnLRq0VCYq+8ypQ/NDiAKYJil2Z5Y
O0t8TtBR7D+3PZkP21OxGBIrfmP2CqBGLflCoPMy69rUbj6LKzHUnMrwSIRKilk2
8TIzC0fxRVzuB4gKrjPQJZ3so+brw9wuUkdmwqR2mU1Asr7X1CFajyE8AYVRylyN
NqjkFsu2bMq7q63tGhPJPCD64u+ke+ooRwHKZ58Y+TwSYEyE7fftvimrqccd5FQa
/84I7dqvWsSIVFfRq4awH+8Q69FAILqjEZYHitRgkOzAB9wwbJns1w2z8/TUfFc3
wEOl9fz+cmqdDH5oxlkXTrzVe/9XbshatARBabeGPE5A3IGoxlAm3/8ij786vs2D
rYV10ZfTNiSUCtx6pFbNoLIO9U2GwzpW28Se2wBtiPqRAomZ1wfGrbJk80xLylMC
4T+gMQxomnmC3cQ6x/2NW7ir61Gg5VN66xYltJgroNZFkg4K4a65+l8wngQU9w9O
XDPuAM4GbRIczBELQ6KZehFZmHi8IMTyrn0dcYYD+pCSnIOU8hr20331+wVuGnQl
BAe06tGrtPGi8ndOA3yhDHofQgAqR9KVgbcL0uZDuU7QhZrG9wq66ow/Yb5HVy0R
NCLgeXVohM0XN98GN8cCghX04ZGhFcpV8NdaoY3jMLbDGyr8AC/2UPgsP0GCn4fr
RnkJqGASdFPgn33YZyiXouaUnHRL49+MsPoO/+GNMY2MqlYDehK4H3nRsEsfISRL
0ZrCvq/zQOmUN4lYhi9BCKqDPJTHeQbKVBEC9ZfdkDddMY/FRYDlI4rjwXJc1I+o
5DeXC+M+UPw/YSJCQFAYG15vI6nfPOWk8FULRwTmAZXM+lJZPnXqc9ntaXYq55NG
Cs9dt4radpy37Y1IZsugn926WjWCZ4E1nFdml66zmdI5oAfZI4aOPm3ivDg8lhnH
tgZ19LdIcNLX+gNQLfsmmc3RxTmKh08ZPbPJLaWzQMgN31CWvgw+MESjrT0mWvY5
f7AsiSve1dZBYUmJCnqrJFMNX13bDHmORhZnMxqKxoW1I2KI8f3eEfpGrLA9lpI0
pmrX/slyGYmchLPYLPDCpR0ciwR/gRPHuMX+DCqUle01L6XtneaCu6bPqLlXper1
WLXIf3bgmhiEoYlPUSmd9FWcXwvoDV5uw3SqnBqjmAdE5D+T+6EyOo2Gg7oJOyh2
s4LrLGEqwXDVCVwAAGiz0xIV+762v1egTxGDqX6zK3vvj4pU3ZpYcEjTpY5CHeUO
ur1400l61jnwIwA0M/bsfL2c9oPhQB70Jgoeyi6aF0Gc4yZCIKCNCmcDtg6P16EW
6x6XzaEVZQzr0NT5AKdwRtrs93ejjAGwSvLtVLtyFUxv7L/QlAB7919chyCSEPs6
+Qr6qCutiFpaTjTCmkQY2LZ5+WKgYLERgbQiYY0t8IA+Q8Bp3sH/9S67CbJE1PQv
b6dIk4e9YvSp/Tk+9Rn7gLB8Cpj8ZE8y7lcyUGoEf3GOcwq086RWub6neCma4K1Y
LRMCxsaYuLCOrr/qsh9z0YajIMyay3EqEmRZCsYlFxwzFQeJqojLGcGIMiRBvDPZ
idakw4h8/U6zIGdQfy+o9X1lJh+DmJRPVlkDXeeFubcG+L2ilKNszxfADVT8ag1w
p48USOZqnHOX+84aFlD6veZu9Bw7PZb8L4Um2rfHwkzgTwBluWp4nCXjXCbyL17z
S7ZAwZXYuBIqoja/egI9yvFhAhwfJbzc5oPzL06dqSnDt4ilMRh2BzoqlArKcrv9
pP70KrftgBlyXt0TLo2djrB7yWtVN576ye1ykPzOrJY65KS534x8QS+y16f1oT/v
tpRLlB8sjomRvYvQ/uDStpl07aIbW0kz0KvqrM3ocqpAGCY02/0hvMIvIw76AHXV
sv+f01L6dX/siVULoQXqwQQYwkrUp9h1hHibB2n1oum8cOEMaE7XX2vJEgD2mxeg
I8ZWdYYf3ow/tiK+DSd8qKiFPVpf/BFZrlqZj+qNs3//jsiuDLonni0K8a6LJZEX
LAFfECTr2kfT/QprVr2ILZHWkaM8R6rmhnPUkTS7qzeFcZ4AMG5sNu2d6QGXtyhP
bXg44FakJdl420Hb4SH2o4xue02X5zLegpOyNPD2FsvJBEVKNSgbtp1W8L5ANazd
P7L9CdjWR8ZE1u7VDDLxmfB/ggukjvgI9QO6ScBEZ7DPNj6lKuGuRDzfJdxyDD8y
CPT4kawB/2tcOWYd5w/enzNe5RcKxO2/HL9vLYTBK4EHkSaejM32r0HE8suaWgX0
2FuBd5oSY7+cu5JmIA0zjbJjfoEFYAvYr8gXJYK/7bw3ooqZTsuw9olYu/KdvQdZ
jpr2J2Imt/BS+AdtIzwSW9kqt54N9Mb5onr9Hfw2DBOlDgO1xpH8GOXFQs+8gJbS
sVbHFziutjOHYVKdndrwtxg41G1jRgNe0ZUkUsoCcX/UqFmpi48JkRbkR+MLBH7V
acFXPIcZRGYs8gHeRe7aBwIeXLZJ0RbPXYEG9dadirqbW9FWbjJeCqfFrOfI29jv
FcVzj3pW09QutAvb9kcqIBRLFyupCbR5H5lHuxLTOk8tZmajeOFF75Otdh79WQw0
uinqLDFXcebrgrwcA+oVS3YA2TCb++n5PZmpKS4+xTVyCfvJxzRyaSybqdKHZ2Eo
ske0x3JKJr8ieSJRMucCHSBoFyE0yUePFdN9pTZ6lwThGBCX9o8Gn1zQLa9xwUxE
+9xpuBfrMlMHOmPKVEQzfJJiPHvImw7ar6T1f73g51HZjvJQce30a12718bPUWVh
YTWNvRUEvwdDVUUB0c6T1iJRd+EUasm5fgQFN2vg0e1b1Lp9leCVfcuUkMeiOcW5
oU57OYi/Y2eoPzRmYxdcPis9MGh2Elumci2AnH7vg66E6jfAEHeHx6N6MieNpXIb
ouxa0WVmoED0/LToegF78aEmZrRfd9tYzcJN/8odgISVXUJWviH1sj4oKpbgO+0x
nlDlHpztkcdnGocRkH3zrqYX71NgTQs34ZoKy4qBuzwbje1yWiC4dJuepDpPOR5l
CHn9W4R6yt9DDrML/08/8WBgd9zpp0Nl8r6fCt+L+Eh7nLTC5dEjcZ95dsfWEX/C
WqjJwrdsS2eVASsDfG0pB6hxT+0Wo0TqzQOIAJAjsYRd4AJEGaFLQol/haf8bRUU
E8L6J+Qk/rzGQWAKw3Cym3rtaepVt0VVlLNZjVrlvkWv4iqYUtQw0+GtikNb7X7L
B0zfXFOPWZd3aQ8DzAReEh0fcca4M1GDQ+jxPM35BzPn02c1BbQJ+GV8YOHwG2+q
orrfr5Ilt0A9uV5Il6YrrY6lLyFmF5dJwBuUGIN9A3qF/JL+PzTP3jfZoC6u6jOU
4DeDsGiHl99edZKxALcHR/kqPREZw+KkNQEiS4VVZmtZKfoMrUwfFOUOEzKQeq3a
Bi8XY9bkv7oEh7XLuGf6B04y4u1kBX/iHPz4f2ofiaYUHpP2jTD+CzlAhsNhaDcB
2kdIEYHnKeDAjjq50cRrY6MXbw7GV9Wu8UyAIdUdPds3vd4l9Phy99in0uQFWKz9
0CkKD8qYWsyNn2Yb72pfp+jYU6V2ocaOiBNV8p/p3xyXnW+juvHUCvQyDWZE50YR
Siey9MeBUjxKDIn9iRciBrjkXgY8Vyx6NIWj+Rj85r9R3AmXZZMwArO80RDWSZkk
1WeyrD+rjuYjmNHDsz1ej0zoF4YaYF7sddhbNKDdSe5rse0TXd0HZ9eohDh8IDmj
MBbhynAZZXo6ZJp3eX+RVjr7xBa3vG5IiKYAUo9TkV1SvLrIy7e8AC5WKPWIwhdx
beINBN91jngzuK0K0cp24t1qIf37UOPEc0Trvi7HzLHDtZMP9egSiL1Urd2G/VhP
bZQp0dD4Rsw33q+CPxV7Xp0z7KBNrizvJeEGIU1FRacrtOvjCTAJyfq/cDb7iPIJ
qL8gKAiebrkiS4Yl7TvhZPmYJWkHUX6Nuant1b1dDgxMaH8yGBzfVbaE1toH4eY7
1uMmnW0+oU5xYaqKYL9zsCSlsrIdUlE3anKZww/RGN29StFekf1k//cWXbVAoav4
ZDudFk2/RbF54zaxLO6RGJIrmGmJr5WZNZtz1kQWbtYwRDcif9ZFDseozjD0fqUg
SASDMTeOVAAuMcchRWyAOvfR3Yw8eQCAx4ua4QgShx3bgGqpf51VZ57eIkhUJwzO
0o13n06y3q2mTgfX0tmWxRuwAIB0N38mBNBZBqsqhLF10l9eMqgCnLTplf9N7oLk
DeAO0O+5hq3FnX0OLz+E9opB0xW9I181IPlGyP18+APr3bP9g6h6r1EP5BcLIVry
opEIStvYb0H8s7HE14P6H6/4+ZuVoZX9ZI2elC62DZb1OSftyi1iH62U8rKLRQ8w
h9wRwQShwlG9WIsdizfimfDL7gOOP/DW/BA873TXFvrOfHmCE/8buOHxwrIm6mFp
swcgQYIvF90evUaNV7pSchf0N61PINhSgO+TCBBDh3YVSaFuS8wY1fN9y7+c3O/a
SFUcKa93rWCrsc/NoT3oWJNbRZWPsZk4Ui4qAKZgeAxMiYR/UCoOll5vBXR4Y6k2
cgk4Kr1A7m/3XnVMOYvT06//oCNskjVjxgOAamm2xWKs1JFw2d0DRCUkNxGhNBUR
TwpC1ism0AdtzZ8oGIWvnlLE226LIiXs5rdZ7FiW3g9A1xYDLBlDEyxTW+T5R1oQ
car5xGVkJQomNBiZ7/ABy8kB9vnS+WuBoI4HP50Q+Hbzxclq+whRhKocgJP8lP2o
xUQZLrsw6HL6sHnLvY53g/6XJYqZUczwnkDl5xiWugW47k7IiNONZn/NMuL3aS32
4/9RgozFCw7isQqsJfG4MhCJGl+5jWjUX187InKcRO3CnZFJyRip1oTklWkFu+h4
EeKpR8uxbIQrjlpdSTUfPVvivpDmSbZfnrJ1m6P4frdmehkGvgSZrlYz+U4/+IgU
lEk15sAIx0T4a5QUe3wSGW2hri8FhPYpWdx7r+jV9CqXpXmx6QrwULJQefzMx6Gf
jft64Vl0uiRJOgtyqY8yctGpyapmC5TvwYGMV37TaA1kG6WKZDRXHjV5S4145gLY
vS3mxQWIKmS8q0tHmuhQ2GPTzrJtB7kaE6PnsBaUAEV5+IUuCgEoQRspblw5dGqK
Y4+uI8QXHX/ka9wENDloYnbJW77iCNXJQ2wsR0aSDtvN2wYs5SONOlA/pzgK/v+6
vCYsU6OINBq1uuPStR/2y6DPWFzGVj0sneKOD+td+WS8kp+RGpzgGIr4K9pxz11M
t2BSQtKTquNwQl89e5w4fMvoFtwT8ecvzA6a5m0MSl1NKGEjZZpXF4bEcd+S31j2
yIgs6M2i2dVPVV9dF9bIRxVon0iXXBhfVBG7dr9x+I894aZR3g1CTkJkXTDSn8rY
1szhQsXUhtJXl0pzCp4KUJ4W30fDRAW2xGOFr60SS4/dPOmNW8pctLnoEF8a65DA
hQB9w3zxg4V21VHK5wMJtjlK1buEAAksXYOurLI6cxoxKX+k2k1AhmH4jG8XDXrt
Vcw7pfDL46TfHyVqwlt7fa9RZNNng8XZH4lz4/ZXZOo4MbBH+t++gSdCBROc0ota
GQgXopjJhK3nTGm0+8SI1kbOEfTEZXJdX0UdCr7LWXbowchp5KrPY493+A0deD9p
5jbtziPOM3CiaaLfHOgZwUA0v6zyV5t85A3LWTGEUXNA/o9ybT8nKkaOg6DkRyeL
lPM3dtXCLjyVOS3ZfqSf6YgRTXH8QHMPEaeoEQjkxk2TfX38VrIfbi/Az4jse97o
KxZ2sgdhTN/QNAZkjVCbMaXTvEKuozNE1LbqK9nI78kKoJeUXxweDQOiHoS2/FaZ
Rgoh3ByqZHa4PEAchYILQva3kanILrnJEa3hFrO5stnFAmyQZXMJkzsMScnmeqSC
iZ6eC/G3xP08pX6jzRAhc+HaRHNm3i+VK4EgVCFMMDYAb/PrHmf0h1uQJf8O1Rxu
/nlfQ/8/lnSB2W85scO/VyABvWfEpgcUiEWdmVQphp6tY/0yNilyOG7aJFy7ol4A
BGHl+vu7ChrEVU98aUGqJr4tq0782ek1NDkD6qHbJu2r82E5SuM2EHE2uH/Nu/W+
//g0TY0sVj9Yv998X9grearp+wTQOj7kKW4+xDKlVLNs0GEfXsazFywmw9FuQs0X
1/Lj249acwwYwzZUm+xKCLRfRkNmtMJhB3GJAo0Vhphc7zw7txyIeX+aXhNT4ww/
JoGjaCUFUzlJZSqAQ4in+FhmnNHo0bDUkWKmsLWFOAynMbMRtd3cSzmW2ko80MFp
afzvz1GnMuCooVJL16aBM52/uINYWDCAKiW2etCYlgob3+RsgzWVaVYS7a16d0SB
q50rqIthFXzO9FerjscFryQYF2yLN4mE4fP34Hx0rjXhb8D6LoEY3J7hpcN3JzS2
6ufh2qb8lL3HlFC9u5VISbTaMp3PPgUN84Yh1eudWVGfH7yxGysBMBBI+/B/I+Eq
bO6ce96Vneu8X9qMM9eTCx4eaB3IMJ4sFBtFIEhU+EAo6TiC7Vhh/gN5KSlluo/Q
4/6mxPSwlLyM+mSxGSvhaAnuuceNB8cKbxIoFpBuyigGlUL+n1fx8lsY+UOL8ysK
W2tUlgWmAndW+dF8j3I66HpxW+aZp9E8zpvuDUkRqYqj9KYSuVnEnWJH0ceOup+L
YZjAOgjAQMabtWJOXOsl/9buX3xSTKHDwIDTeBktR590TDOVqn+DmITXemK4Czb4
MOq/4JiOKWxo4doJ2IUVLrzl9m57WuXsoWVdp4EwPVGFSECcC+3aTWqcVbgn8FMP
wSwMaY8r2VWkgCwy0Bin5NJ+4d0t1RywghuzyK/QrcmRVdc8WJ/zE1oBZLLhO9Wx
c6WUakWDf5is8h9W5ogZJibyo1p3NuCx0CqxFNceTPDo1gr6V3lvIAeHIyKpi7Et
dHqwFGS+7dcMjF1YlLvpDBfLs9fVnSa6Jb2Asyv3uXSqhQvv1X/qshT4n1d74I3c
P21VOTxXneTUMI0KDrAHbJRvs/D8uUEg+xVC1DIGpzmnQua2sqL2zu7qulA/jy51
tmcrN4V8t995F++vX6oM61sH7hIuIU1Qa9dfP3vtsnNjlh3BvhFtPvTBFF5hfv8v
xIFOtMNCyXS2jLL3eBwP4VhtVPOCQFPV7P2tsNJq/ih1aNhHnlMsl/QTEt1Ynk0o
Ilvpgv2hNEgnXY0tlWw8ekrOPUIRJZgf5NkaXJ0mU4ukG+i55dkP8TSiDgnHguLH
YRuCu5+dE0Wgtm8qfvHFfqR5zQWhhMQVE+6FsuAnNi4iygADphPb/b9QENTztxlC
C1h86LHD75aAuyKaq367QUezvtbzOpWI28pmqzfh/mY0TaPUoEua72GxfCk4r0sV
LOOa5Xx6ySpWwwtCovgdkENUxraL8hUGCmlqKilWzD6+lsaOYPLOGYcjihQx4uIo
ptbi8FhLkCNEzNsth9mtYNJIqUfDtW/hmTEDBzK3LDOzywTfqF81In+EIp5sMQ/N
XuyYmKV/tSQb8smHQZs/dsPyvutHMQpeKNm1208nQDYYCfCIans+cBzQ+bJVQ3pX
Bd/D3RAZ8D/FGn4Q4Gy5G4LMLMTwirOJHJJscc8F7zBTOQY4bMD9rEGH9RVs3Kmz
d0egxa5K53HMTNfFCv5cSF7wZr1FOniyihIUQqmsmCCeWr/iaz3sE8yyGdaXenB0
SYyTCM5SWWr0mL/S5nHYEYHRWwLT8ccJM97WoVWkYNJeXcI83dafQnEWwKlrWPHB
jZGm96c9izc/GsYlZg5DVfufyCy6Y0HhFyd/Rr+y4U/2bDVkN9jY/Bx4bYprIc4I
d1KhYkEO5UUNZjITApAZ1wem2+tZiWxX6Teaqev5AN2/XeYI2Pe4PCjvHrCbGMse
0wGabXGkfmgS4kI4bIWJ/jfgMDQq66MLKPDz0kX7BBmDKDF5B7XHjZTtnmHzIfoZ
3zRwZy4OA2927GAu5b7msgao6ngurGjZ2YyAQfdqf2xtdK9OUZXcHG6RYE47+IlD
b83uXkUe/KXBiOhV47fi8Hipv4dEq/TEgvfrVuwASxYZS760C4G2nCCEj42H2PAF
4Ni7xlh8WNpv5b9522/rhrMhJZ4pZHJThLo8nxIpu8+LifoR5AUiyD0i7yMNA+FB
OVAxE2GpGWvWoTf9MPp+nwsHPuLfq2LOQAQT82DOb0ipj/VQXb/59iSP3oL5Snbi
lmS1bW34iKrIYqvtWeuYKC3D8t542SfkkPyTkg5XI3yCfcNQ4JIucs4fqQ5d8eqo
OE4YPbtqa9kyI5N3cKMDQOlk2hBjShCttVdpXAaQvcmid7Ew9gjvBdsSD8gt1/EC
q6YBdnAaZ3V/nzVW+m+TR8PzkTicof2BwGfRNq1chJdIoKmDH8nVDbSpdzBXJbl3
nCNkLL153hLucKXrycGPupy4sb2nx/kUVmNLq913goDugNDjO1c63G+M8Nq0BUah
efRjp6iwg83+2Z/TmjYdLOJUIRs5OAvVp2hwquP3YWOH/XQnWth4idZXj3R4KWnl
xI8SCs/x2RKsqjb22Jzni7WPQLW0DHsxXixZENrSCDqkzJcIBcCe39thwx6FUtWZ
gA8OjkmR4wvI3Ibnkl+MU+jlEV1GZRGEUn0WArNhgkHJ5PnOnOi026tnUsl6JeIc
6nmpo/bmwvB5KeFLQAGL6Kcs5SuFy0q2RznphOzl1WBcLH/KEOSM1cfRhG4B4+IM
2nLHV+r7o0u5tWgc+lyt1JN0fRPMNXEWJ1KT1lGcuhIrEs63RrA3YlyDmbmb8oiZ
OH3X7TeNK2T33cWQ8JGQ387n4KRz0RqAN8cklLm71fzZFbDT8riTTtMC1Mx5RawF
/TuophPRYoxFxaSfZeAIImZLSYt9frldPsK8WHEbw5srrLY2HFOWWZ70OSFVFCEu
Rnx6y6Onk70yTDvQ8dOUETBbF1JZYKW5RHy+ZXVWlMxHi+x7xVRhs3VVM0zpeMN2
N89200LMIejVg/g3NKMx5y9B2HIz10D4ZPamywGHAAW88ktxVDqq5zgnyf/Cc8C7
THatMxVA1uJ5JSRokiad5jwuogA3PaXDYFtemo9AKVHjL4f5ULl7TWcWJKum7B36
tNsIRY+uWJ7E70ArzXxJXCJfYpypYsHrAN0yzrNlvu/WrBGmZgsS/FAgQ0G4mi4B
p9lMjmU/A9KNn4zBN1+hOJ9JnCL9273fJezrJbocapnheVI7szU6RR7Jhy+yXIVC
udQIeaYV26iq97MTh+6vHS+toLaAg9R2Xrj1f/H3hZtW2lEJ5MOrvhS2xeYYKp3w
hKFm4o97G7PIyOB5n0JSWGzUiMbwNILlQ+WGQJx4ZG7XW3AbZvGmDWqeSu6mqmf3
`pragma protect end_protected